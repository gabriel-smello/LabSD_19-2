library IEEE;
use IEEE.std_logic_1164.all;

entity exp8visto2 is
    port( clock : in std_logic;
          reset : in std_logic;
          T60 : out std_logic;
          T20 : out std_logic;
          T6 : out std_logic;
          T5 : out std_logic;
          num7seg : out std_logic_vector(7 downto 0);
          displays : out std_logic_vector(3 downto 0));
end exp8visto2;

architecture exp8visto2_arch of exp8visto2 is
    --inserir sinais e componentes aqui
begin 

    --inserir implemnetação aqui

end exp8visto2_arch;