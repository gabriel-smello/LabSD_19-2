-- Somador de 4 bits usando apenas somadores completos.
-- Utilizar visto 1 do experimento 2 como "component".
-- Dois vetores  A e B com 4 bits de entrada.
-- Um vetor S com 5 bits de saida.
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;

entity somador_golden is
    port(a, B: in S);
end somador4; 

architecture somador4_arch of somador4 is
begin
    

    
end somador4_arch;
