library IEEE;
use IEEE.std_logic_1164.all;

entity exp8visto3 is
    port( clock : in std_logic;
          ligadesliga : in std_logic;
          sensorA : out std_logic;
          sensorB : out std_logic;
          num7seg : out std_logic_vector(7 downto 0);
          displays : out std_logic_vector(3 downto 0));
end exp8visto3;

architecture exp8visto3_arch of exp8visto3 is
    --inserir sinais e componentes aqui
begin 

    --inserir implemnetação aqui

end exp8visto3_arch;